--
-- Copyright 2017 Gary Preston <gary@mups.co.uk>
-- All rights reserved
--
-- Redistribution and use in source and synthesized forms, with or without
-- modification, are permitted provided that the following conditions are met:
--
-- Redistributions of source code must retain the above copyright notice,
-- this list of conditions and the following disclaimer.
--
-- Redistributions in synthesized form must reproduce the above copyright
-- notice, this list of conditions and the following disclaimer in the
-- documentation and/or other materials provided with the distribution.
--
-- Neither the name of the author nor the names of other contributors may
-- be used to endorse or promote products derived from this software without
-- specific prior written permission.
--
-- License is granted for non-commercial use only.  A fee may not be charged
-- for redistributions as source code or in synthesized/hardware form without
-- specific prior written permission.
--
-- THIS CODE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
-- AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR
-- PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE AUTHOR OR CONTRIBUTORS BE
-- LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR
-- CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF
-- SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS
-- INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN
-- CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE
-- POSSIBILITY OF SUCH DAMAGE.
--
-- You are responsible for any legal issues arising from your use of this code.
--

-- Interface Frequency based ULA cassette pins with SD Card based 
-- files using Generic FileIO.

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

use work.Replay_Pack.all;

entity Virtual_Cassette_FileIO is
  port (
    -- Clocks (32MHz sys with 1:4 enable)
    i_clk                : in bit1;
    i_ena                : in bit1;
    i_rst                : in bit1;

    -- FileIO channel
    i_fch_cfg            : in  r_Cfg_fileio;
    i_fch_to_core        : in  r_Fileio_to_core;
    o_fch_fm_core        : out r_Fileio_fm_core;

    -- Tape Controls
    i_motor              : in bit1;
    i_play               : in bit1;
    i_rec                : in bit1;
    i_ffwd               : in bit1;
    i_rwnd               : in bit1;

    -- Pulse based cassette i/o (0 = 1200Hz and 1 = 2400Hz)
    i_cas_to_fch         : in bit1;
    o_cas_fm_fch         : out bit1
  );
end;

architecture RTL of Virtual_Cassette_FileIO is
  signal data : word(7 downto 0);
  signal dummy_addr : integer range 5000 downto 0 := 0;


begin

  -- Temp disabled until file io hooked up
  o_fch_fm_core <= Z_Fileio_fm_core;

  -- File IO only handles 0 or 1 states where as tape had pulses of 0's
  -- pulses of 1's and then gaps with level 0. Gaps will end up generating
  -- pulses of 0's with the current setup. Although this should hopefully
  -- not cause too big a problem as the first run of 0's will cause the
  -- stop bit check to fail and a return to looking for a high tone.
  -- There will be a single byte that generates a RX full interrupt however.
  
  -- For initial testing return an incrementing counter for each byte
  -- to verify the ULA's side of the loading works, before complicating
  -- with FileIO.

  -- Assumes start/stop bits are baked into the stream already.
  p_dummy_read : process(i_clk, i_ena, i_rst)
    variable cnt : integer := 0;
    variable cur_bit : integer range 7 downto 0;    
  begin
    if (i_rst = '1') then
      cnt := 0;
      dummy_addr <= 0;
      cur_bit := 7;
    elsif rising_edge(i_clk) then
      -- TODO: check inserted etc

      -- temporary position reset to ease testing
      if (i_play = '0' or i_motor = '0') then
        dummy_addr <= 0;
        cur_bit := 7;
        cnt := 0;
      end if;

      -- Hacky test to load part of a acorn tape which has been converted
      -- from uef to a bitstream including start/stop bits and then pasted
      -- into a giant case.
      if (i_ena = '1') and (i_play = '1') and (i_motor = '1') then
        if cnt = 0 then
          if cur_bit = 7 then
            cur_bit := 0;
          else            
            cur_bit := cur_bit + 1;
          end if;

          -- i_ena @8MHz
          cnt := 6666;
        end if;

        cnt := cnt - 1;

        -- Ready new byte by next clock
        if cnt = 0 and cur_bit = 7 then
          dummy_addr <= dummy_addr + 1;
        end if;
        
      end if;      

      o_cas_fm_fch <= '0';
      -- Pulse generation: 2400Hz = 0, 2x1200Hz = 1
      if (data(7-cur_bit) = '1' and cnt > 1666 and cnt < 3333) or
        (data(7-cur_bit) = '1' and cnt > 4999) or
        (data(7-cur_bit) = '0' and cnt > 3333) then
          o_cas_fm_fch <= '1';
      end if;
    end if;

  end process;

  p_data : process(i_clk, i_ena, i_rst)
  begin
    
    if rising_edge(i_clk) then
      data <= (others => '0');

      case dummy_addr is
        when 0 => data <= "11111111";
        when 1 => data <= "11111111";
        when 2 => data <= "11111111";      
        when 3 => data <= "11111111";
        when 4 => data <= "11111111";
        when 5 => data <= "11111111";
        when 6 => data <= "11111111";
        when 7 => data <= "11111111";
        when 8 => data <= "11111111";
        when 9 => data <= "11111111";
        when 10 => data <= "11111111";
        when 11 => data <= "11111111";
        when 12 => data <= "11111111";
        when 13 => data <= "11111111";
        when 14 => data <= "11111111";
        when 15 => data <= "11111111";
        when 16 => data <= "11111111";
        when 17 => data <= "11111111";
        when 18 => data <= "11111111";
        when 19 => data <= "11111111";
        when 20 => data <= "11111111";
        when 21 => data <= "11111111";
        when 22 => data <= "11111111";
        when 23 => data <= "11111111";
        when 24 => data <= "11111111";
        when 25 => data <= "11111111";
        when 26 => data <= "11111111";
        when 27 => data <= "11111111";
        when 28 => data <= "11111111";
        when 29 => data <= "11111111";
        when 30 => data <= "11111111";
        when 31 => data <= "11111111";
        when 32 => data <= "11111111";
        when 33 => data <= "11111111";
        when 34 => data <= "11111111";
        when 35 => data <= "11111111";
        when 36 => data <= "11111111";
        when 37 => data <= "11111111";
        when 38 => data <= "11111111";
        when 39 => data <= "11111111";
        when 40 => data <= "11111111";
        when 41 => data <= "11111111";
        when 42 => data <= "11111111";
        when 43 => data <= "11111111";
        when 44 => data <= "11111111";
        when 45 => data <= "11111111";
        when 46 => data <= "11111111";
        when 47 => data <= "11111111";
        when 48 => data <= "11111111";
        when 49 => data <= "11111111";
        when 50 => data <= "11111111";
        when 51 => data <= "11111111";
        when 52 => data <= "11111111";
        when 53 => data <= "11111111";
        when 54 => data <= "11111111";
        when 55 => data <= "11111111";
        when 56 => data <= "11111111";
        when 57 => data <= "11111111";
        when 58 => data <= "11111111";
        when 59 => data <= "11111111";
        when 60 => data <= "11111111";
        when 61 => data <= "11111111";
        when 62 => data <= "11111111";
        when 63 => data <= "11111111";
        when 64 => data <= "11111111";
        when 65 => data <= "11111111";
        when 66 => data <= "11111111";
        when 67 => data <= "11111111";
        when 68 => data <= "11111111";
        when 69 => data <= "11111111";
        when 70 => data <= "11111111";
        when 71 => data <= "11111111";
        when 72 => data <= "11111111";
        when 73 => data <= "11111111";
        when 74 => data <= "11111111";
        when 75 => data <= "11111111";
        when 76 => data <= "11111111";
        when 77 => data <= "11111111";
        when 78 => data <= "11111111";
        when 79 => data <= "11111111";
        when 80 => data <= "11111111";
        when 81 => data <= "11111111";
        when 82 => data <= "11111111";
        when 83 => data <= "11111111";
        when 84 => data <= "11111111";
        when 85 => data <= "11111111";
        when 86 => data <= "11111111";
        when 87 => data <= "11111111";
        when 88 => data <= "11111111";
        when 89 => data <= "11111111";
        when 90 => data <= "11111111";
        when 91 => data <= "11111111";
        when 92 => data <= "11111111";
        when 93 => data <= "11111111";
        when 94 => data <= "11111111";
        when 95 => data <= "11111111";
        when 96 => data <= "11111111";
        when 97 => data <= "11111111";
        when 98 => data <= "11111111";
        when 99 => data <= "11111111";
        when 100 => data <= "11111111";
        when 101 => data <= "11111111";
        when 102 => data <= "11111111";
        when 103 => data <= "11111111";
        when 104 => data <= "11111111";
        when 105 => data <= "11111111";
        when 106 => data <= "11111111";
        when 107 => data <= "11111111";
        when 108 => data <= "11111111";
        when 109 => data <= "11111111";
        when 110 => data <= "11111111";
        when 111 => data <= "11111111";
        when 112 => data <= "11111111";
        when 113 => data <= "11111111";
        when 114 => data <= "11111111";
        when 115 => data <= "11111111";
        when 116 => data <= "11111111";
        when 117 => data <= "11111111";
        when 118 => data <= "11111111";
        when 119 => data <= "11111111";
        when 120 => data <= "11111111";
        when 121 => data <= "11111111";
        when 122 => data <= "11111111";
        when 123 => data <= "11111111";
        when 124 => data <= "11111111";
        when 125 => data <= "11111111";
        when 126 => data <= "11111111";
        when 127 => data <= "11111111";
        when 128 => data <= "11111111";
        when 129 => data <= "11111111";
        when 130 => data <= "11111111";
        when 131 => data <= "11111111";
        when 132 => data <= "11111111";
        when 133 => data <= "11111111";
        when 134 => data <= "11111111";
        when 135 => data <= "11111111";
        when 136 => data <= "11111111";
        when 137 => data <= "11111111";
        when 138 => data <= "11111111";
        when 139 => data <= "11111111";
        when 140 => data <= "11111111";
        when 141 => data <= "11111111";
        when 142 => data <= "11111111";
        when 143 => data <= "11111111";
        when 144 => data <= "11111111";
        when 145 => data <= "11111111";
        when 146 => data <= "11111111";
        when 147 => data <= "11111111";
        when 148 => data <= "11111111";
        when 149 => data <= "11111111";
        when 150 => data <= "11111111";
        when 151 => data <= "11111111";
        when 152 => data <= "11111111";
        when 153 => data <= "11111111";
        when 154 => data <= "11111111";
        when 155 => data <= "11111111";
        when 156 => data <= "11111111";
        when 157 => data <= "11111111";
        when 158 => data <= "11111111";
        when 159 => data <= "11111111";
        when 160 => data <= "11111111";
        when 161 => data <= "11111111";
        when 162 => data <= "11111111";
        when 163 => data <= "11111111";
        when 164 => data <= "11111111";
        when 165 => data <= "11111111";
        when 166 => data <= "11111111";
        when 167 => data <= "11111111";
        when 168 => data <= "11111111";
        when 169 => data <= "11111111";
        when 170 => data <= "11111111";
        when 171 => data <= "11111111";
        when 172 => data <= "11111111";
        when 173 => data <= "11111111";
        when 174 => data <= "11111111";
        when 175 => data <= "11111111";
        when 176 => data <= "11111111";
        when 177 => data <= "11111111";
        when 178 => data <= "11111111";
        when 179 => data <= "11111111";
        when 180 => data <= "11111111";
        when 181 => data <= "11111111";
        when 182 => data <= "11111111";
        when 183 => data <= "11111111";
        when 184 => data <= "11111111";
        when 185 => data <= "11111111";
        when 186 => data <= "11111111";
        when 187 => data <= "11111111";
        when 188 => data <= "11111111";
        when 189 => data <= "11111111";
        when 190 => data <= "11111111";
        when 191 => data <= "11111111";
        when 192 => data <= "11111111";
        when 193 => data <= "11111111";
        when 194 => data <= "11111111";
        when 195 => data <= "11111111";
        when 196 => data <= "11111111";
        when 197 => data <= "11111111";
        when 198 => data <= "11111111";
        when 199 => data <= "11111111";
        when 200 => data <= "11111111";
        when 201 => data <= "11111111";
        when 202 => data <= "11111111";
        when 203 => data <= "11111111";
        when 204 => data <= "11111111";
        when 205 => data <= "11111111";
        when 206 => data <= "11111111";
        when 207 => data <= "11111111";
        when 208 => data <= "11111111";
        when 209 => data <= "11111111";
        when 210 => data <= "11111111";
        when 211 => data <= "11111111";
        when 212 => data <= "11111111";
        when 213 => data <= "11111111";
        when 214 => data <= "11111111";
        when 215 => data <= "11111111";
        when 216 => data <= "11111111";
        when 217 => data <= "11111111";
        when 218 => data <= "11111111";
        when 219 => data <= "11111111";
        when 220 => data <= "11111111";
        when 221 => data <= "11111111";
        when 222 => data <= "11111111";
        when 223 => data <= "11111111";
        when 224 => data <= "11111111";
        when 225 => data <= "11000111";
        when 226 => data <= "01111111";
        when 227 => data <= "11111111";
        when 228 => data <= "11111111";
        when 229 => data <= "11111111";
        when 230 => data <= "11111111";
        when 231 => data <= "11111111";
        when 232 => data <= "11111111";
        when 233 => data <= "11111111";
        when 234 => data <= "11111111";
        when 235 => data <= "11111111";
        when 236 => data <= "11111111";
        when 237 => data <= "11111111";
        when 238 => data <= "11111111";
        when 239 => data <= "11111111";
        when 240 => data <= "11111111";
        when 241 => data <= "11111111";
        when 242 => data <= "11111111";
        when 243 => data <= "11111111";
        when 244 => data <= "11111111";
        when 245 => data <= "11111111";
        when 246 => data <= "11111111";
        when 247 => data <= "11111111";
        when 248 => data <= "11111111";
        when 249 => data <= "11111111";
        when 250 => data <= "11111111";
        when 251 => data <= "11111111";
        when 252 => data <= "11111111";
        when 253 => data <= "11111111";
        when 254 => data <= "11111111";
        when 255 => data <= "11111111";
        when 256 => data <= "11111111";
        when 257 => data <= "11111111";
        when 258 => data <= "11111111";
        when 259 => data <= "11111111";
        when 260 => data <= "11111111";
        when 261 => data <= "11111111";
        when 262 => data <= "11111111";
        when 263 => data <= "11111111";
        when 264 => data <= "11111111";
        when 265 => data <= "11111111";
        when 266 => data <= "11111111";
        when 267 => data <= "11111111";
        when 268 => data <= "11111111";
        when 269 => data <= "11111111";
        when 270 => data <= "11111111";
        when 271 => data <= "11111111";
        when 272 => data <= "11111111";
        when 273 => data <= "11111111";
        when 274 => data <= "11111111";
        when 275 => data <= "11111111";
        when 276 => data <= "11111111";
        when 277 => data <= "11111111";
        when 278 => data <= "11111111";
        when 279 => data <= "11111111";
        when 280 => data <= "11111111";
        when 281 => data <= "11111111";
        when 282 => data <= "11111111";
        when 283 => data <= "11111111";
        when 284 => data <= "11111111";
        when 285 => data <= "11111111";
        when 286 => data <= "11111111";
        when 287 => data <= "11111111";
        when 288 => data <= "11111111";
        when 289 => data <= "11111111";
        when 290 => data <= "11111111";
        when 291 => data <= "11111111";
        when 292 => data <= "11111111";
        when 293 => data <= "11111111";
        when 294 => data <= "11111111";
        when 295 => data <= "11111111";
        when 296 => data <= "11111111";
        when 297 => data <= "11111111";
        when 298 => data <= "11111111";
        when 299 => data <= "11111111";
        when 300 => data <= "11111111";
        when 301 => data <= "11111111";
        when 302 => data <= "11111111";
        when 303 => data <= "11111111";
        when 304 => data <= "11111111";
        when 305 => data <= "11111111";
        when 306 => data <= "11111111";
        when 307 => data <= "11111111";
        when 308 => data <= "11111111";
        when 309 => data <= "11111111";
        when 310 => data <= "11111111";
        when 311 => data <= "11111111";
        when 312 => data <= "11111111";
        when 313 => data <= "11111111";
        when 314 => data <= "11111111";
        when 315 => data <= "11111111";
        when 316 => data <= "11111111";
        when 317 => data <= "11111111";
        when 318 => data <= "11111111";
        when 319 => data <= "11111111";
        when 320 => data <= "11111111";
        when 321 => data <= "11111111";
        when 322 => data <= "11111111";
        when 323 => data <= "11111111";
        when 324 => data <= "11111111";
        when 325 => data <= "11111111";
        when 326 => data <= "11111111";
        when 327 => data <= "11111111";
        when 328 => data <= "11111111";
        when 329 => data <= "11111111";
        when 330 => data <= "11111111";
        when 331 => data <= "11111111";
        when 332 => data <= "11111111";
        when 333 => data <= "11111111";
        when 334 => data <= "11111111";
        when 335 => data <= "11111111";
        when 336 => data <= "11111111";
        when 337 => data <= "11111111";
        when 338 => data <= "11111111";
        when 339 => data <= "11111111";
        when 340 => data <= "11111111";
        when 341 => data <= "11111111";
        when 342 => data <= "11111111";
        when 343 => data <= "11111111";
        when 344 => data <= "11111111";
        when 345 => data <= "11111111";
        when 346 => data <= "11111111";
        when 347 => data <= "11111111";
        when 348 => data <= "11111111";
        when 349 => data <= "11111111";
        when 350 => data <= "11111111";
        when 351 => data <= "11111111";
        when 352 => data <= "11111111";
        when 353 => data <= "11111111";
        when 354 => data <= "11111111";
        when 355 => data <= "11111111";
        when 356 => data <= "11111111";
        when 357 => data <= "11111111";
        when 358 => data <= "11111111";
        when 359 => data <= "11111111";
        when 360 => data <= "11111111";
        when 361 => data <= "11111111";
        when 362 => data <= "11111111";
        when 363 => data <= "11111111";
        when 364 => data <= "11111111";
        when 365 => data <= "11111111";
        when 366 => data <= "11111111";
        when 367 => data <= "11111111";
        when 368 => data <= "11111111";
        when 369 => data <= "11111111";
        when 370 => data <= "11111111";
        when 371 => data <= "11111111";
        when 372 => data <= "11111111";
        when 373 => data <= "11111111";
        when 374 => data <= "11111111";
        when 375 => data <= "11111111";
        when 376 => data <= "11111111";
        when 377 => data <= "11111111";
        when 378 => data <= "11111111";
        when 379 => data <= "11111111";
        when 380 => data <= "11111111";
        when 381 => data <= "11111111";
        when 382 => data <= "11111111";
        when 383 => data <= "11111111";
        when 384 => data <= "11111111";
        when 385 => data <= "11111111";
        when 386 => data <= "11111111";
        when 387 => data <= "11111111";
        when 388 => data <= "11111111";
        when 389 => data <= "11111111";
        when 390 => data <= "11111111";
        when 391 => data <= "11111111";
        when 392 => data <= "11111111";
        when 393 => data <= "11111111";
        when 394 => data <= "11111111";
        when 395 => data <= "11111111";
        when 396 => data <= "11111111";
        when 397 => data <= "11111111";
        when 398 => data <= "11111111";
        when 399 => data <= "11111111";
        when 400 => data <= "11111111";
        when 401 => data <= "11111111";
        when 402 => data <= "11111111";
        when 403 => data <= "11111111";
        when 404 => data <= "11111111";
        when 405 => data <= "11111111";
        when 406 => data <= "11111111";
        when 407 => data <= "11111111";
        when 408 => data <= "11111111";
        when 409 => data <= "11111111";
        when 410 => data <= "11111111";
        when 411 => data <= "11111111";
        when 412 => data <= "11111111";
        when 413 => data <= "11111111";
        when 414 => data <= "11111111";
        when 415 => data <= "11111111";
        when 416 => data <= "11111111";
        when 417 => data <= "11111111";
        when 418 => data <= "11111111";
        when 419 => data <= "11111111";
        when 420 => data <= "11111111";
        when 421 => data <= "11111111";
        when 422 => data <= "11111111";
        when 423 => data <= "11111111";
        when 424 => data <= "11111111";
        when 425 => data <= "11111111";
        when 426 => data <= "11111111";
        when 427 => data <= "11111111";
        when 428 => data <= "11111111";
        when 429 => data <= "11111111";
        when 430 => data <= "11111111";
        when 431 => data <= "11111111";
        when 432 => data <= "11111111";
        when 433 => data <= "11111111";
        when 434 => data <= "11111111";
        when 435 => data <= "11111111";
        when 436 => data <= "11111111";
        when 437 => data <= "11111111";
        when 438 => data <= "11111111";
        when 439 => data <= "11111111";
        when 440 => data <= "11111111";
        when 441 => data <= "11111111";
        when 442 => data <= "11111111";
        when 443 => data <= "11111111";
        when 444 => data <= "11111111";
        when 445 => data <= "11111111";
        when 446 => data <= "11111111";
        when 447 => data <= "11111111";
        when 448 => data <= "11111111";
        when 449 => data <= "11111111";
        when 450 => data <= "11111111";
        when 451 => data <= "11111100";
        when 452 => data <= "10101001";
        when 453 => data <= "01010001";
        when 454 => data <= "01000110";
        when 455 => data <= "01010100";
        when 456 => data <= "10010100";
        when 457 => data <= "01010101";
        when 458 => data <= "01010001";
        when 459 => data <= "01000000";
        when 460 => data <= "00010000";
        when 461 => data <= "00000101";
        when 462 => data <= "00110001";
        when 463 => data <= "01111111";
        when 464 => data <= "11011111";
        when 465 => data <= "11110110";
        when 466 => data <= "00100100";
        when 467 => data <= "00000011";
        when 468 => data <= "01111111";
        when 469 => data <= "11011111";
        when 470 => data <= "11110000";
        when 471 => data <= "00000100";
        when 472 => data <= "00000001";
        when 473 => data <= "01101111";
        when 474 => data <= "11000000";
        when 475 => data <= "00010000";
        when 476 => data <= "00001100";
        when 477 => data <= "00000001";
        when 478 => data <= "00000000";
        when 479 => data <= "01000000";
        when 480 => data <= "00010000";
        when 481 => data <= "00000100";
        when 482 => data <= "01010101";
        when 483 => data <= "00101111";
        when 484 => data <= "01010110";
        when 485 => data <= "00010000";
        when 486 => data <= "00000100";
        when 487 => data <= "10100001";
        when 488 => data <= "00111100";
        when 489 => data <= "01000101";
        when 490 => data <= "11110000";
        when 491 => data <= "00100100";
        when 492 => data <= "00001001";
        when 493 => data <= "00000010";
        when 494 => data <= "01000000";
        when 495 => data <= "10010000";
        when 496 => data <= "00100100";
        when 497 => data <= "00001001";
        when 498 => data <= "00000010";
        when 499 => data <= "01000000";
        when 500 => data <= "10010000";
        when 501 => data <= "00100100";
        when 502 => data <= "11101001";
        when 503 => data <= "00111010";
        when 504 => data <= "01001110";
        when 505 => data <= "10010101";
        when 506 => data <= "00010100";
        when 507 => data <= "00001001";
        when 508 => data <= "00011001";
        when 509 => data <= "01000000";
        when 510 => data <= "10010100";
        when 511 => data <= "10010100";
        when 512 => data <= "00001001";
        when 513 => data <= "00010101";
        when 514 => data <= "01000000";
        when 515 => data <= "10010101";
        when 516 => data <= "00010100";
        when 517 => data <= "11101001";
        when 518 => data <= "00111010";
        when 519 => data <= "01001110";
        when 520 => data <= "10010000";
        when 521 => data <= "00100101";
        when 522 => data <= "01100001";
        when 523 => data <= "00000000";
        when 524 => data <= "01000101";
        when 525 => data <= "00010101";
        when 526 => data <= "00000100";
        when 527 => data <= "00001001";
        when 528 => data <= "01011000";
        when 529 => data <= "01000000";
        when 530 => data <= "00010011";
        when 531 => data <= "11000101";
        when 532 => data <= "00001001";
        when 533 => data <= "00010111";
        when 534 => data <= "11000000";
        when 535 => data <= "10010000";
        when 536 => data <= "00100100";
        when 537 => data <= "00001001";
        when 538 => data <= "00000010";
        when 539 => data <= "01001110";
        when 540 => data <= "10010011";
        when 541 => data <= "10100100";
        when 542 => data <= "11101001";
        when 543 => data <= "01010001";
        when 544 => data <= "01000110";
        when 545 => data <= "11010101";
        when 546 => data <= "00110101";
        when 547 => data <= "10001101";
        when 548 => data <= "00010111";
        when 549 => data <= "01001001";
        when 550 => data <= "11010111";
        when 551 => data <= "10110100";
        when 552 => data <= "11101101";
        when 553 => data <= "00000010";
        when 554 => data <= "01001101";
        when 555 => data <= "01010101";
        when 556 => data <= "00110100";
        when 557 => data <= "10011101";
        when 558 => data <= "01100111";
        when 559 => data <= "01010010";
        when 560 => data <= "11010111";
        when 561 => data <= "10110100";
        when 562 => data <= "11101101";
        when 563 => data <= "00000010";
        when 564 => data <= "01010001";
        when 565 => data <= "10010011";
        when 566 => data <= "10100100";
        when 567 => data <= "11101001";
        when 568 => data <= "00111010";
        when 569 => data <= "01010110";
        when 570 => data <= "00010000";
        when 571 => data <= "00000100";
        when 572 => data <= "00101001";
        when 573 => data <= "01010000";
        when 574 => data <= "01000000";
        when 575 => data <= "10010101";
        when 576 => data <= "10000100";
        when 577 => data <= "00000001";
        when 578 => data <= "00100110";
        when 579 => data <= "01001111";
        when 580 => data <= "00010001";
        when 581 => data <= "01111100";
        when 582 => data <= "00001001";
        when 583 => data <= "00000010";
        when 584 => data <= "01000000";
        when 585 => data <= "10010000";
        when 586 => data <= "00100100";
        when 587 => data <= "00001001";
        when 588 => data <= "00000010";
        when 589 => data <= "01000000";
        when 590 => data <= "10010000";
        when 591 => data <= "00100100";
        when 592 => data <= "00001001";
        when 593 => data <= "00000010";
        when 594 => data <= "01011000";
        when 595 => data <= "01010111";
        when 596 => data <= "10110100";
        when 597 => data <= "00011101";
        when 598 => data <= "01001111";
        when 599 => data <= "01001001";
        when 600 => data <= "11010100";
        when 601 => data <= "10110101";
        when 602 => data <= "11001101";
        when 603 => data <= "00001011";
        when 604 => data <= "01000101";
        when 605 => data <= "11010000";
        when 606 => data <= "00100100";
        when 607 => data <= "00101001";
        when 608 => data <= "01100011";
        when 609 => data <= "01010010";
        when 610 => data <= "10010000";
        when 611 => data <= "00100100";
        when 612 => data <= "00001001";
        when 613 => data <= "01011000";
        when 614 => data <= "01000000";
        when 615 => data <= "00010001";
        when 616 => data <= "11100100";
        when 617 => data <= "10001001";
        when 618 => data <= "00010111";
        when 619 => data <= "11000000";
        when 620 => data <= "10010000";
        when 621 => data <= "00100100";
        when 622 => data <= "00001001";
        when 623 => data <= "00000010";
        when 624 => data <= "01000000";
        when 625 => data <= "10010100";
        when 626 => data <= "00010101";
        when 627 => data <= "10001101";
        when 628 => data <= "01111011";
        when 629 => data <= "01001001";
        when 630 => data <= "11010011";
        when 631 => data <= "10110101";
        when 632 => data <= "10011101";
        when 633 => data <= "01111011";
        when 634 => data <= "01001100";
        when 635 => data <= "11010001";
        when 636 => data <= "01110100";
        when 637 => data <= "00001001";
        when 638 => data <= "00011001";
        when 639 => data <= "01010010";
        when 640 => data <= "11010101";
        when 641 => data <= "10110101";
        when 642 => data <= "00101101";
        when 643 => data <= "00010111";
        when 644 => data <= "01010100";
        when 645 => data <= "11010001";
        when 646 => data <= "00110100";
        when 647 => data <= "00001001";
        when 648 => data <= "01000110";
        when 649 => data <= "01010011";
        when 650 => data <= "10010000";
        when 651 => data <= "11100100";
        when 652 => data <= "01011001";
        when 653 => data <= "00000010";
        when 654 => data <= "01000000";
        when 655 => data <= "10010101";
        when 656 => data <= "10000100";
        when 657 => data <= "00000001";
        when 658 => data <= "00110001";
        when 659 => data <= "01010100";
        when 660 => data <= "00010000";
        when 661 => data <= "00100101";
        when 662 => data <= "01100001";
        when 663 => data <= "00000000";
        when 664 => data <= "01000001";
        when 665 => data <= "01010111";
        when 666 => data <= "10000101";
        when 667 => data <= "10101111";
        when 668 => data <= "01110110";
        when 669 => data <= "01001011";
        when 670 => data <= "10010010";
        when 671 => data <= "10100100";
        when 672 => data <= "11000101";
        when 673 => data <= "00001101";
        when 674 => data <= "01001001";
        when 675 => data <= "10010000";
        when 676 => data <= "01100100";
        when 677 => data <= "00011001";
        when 678 => data <= "00000010";
        when 679 => data <= "01001001";
        when 680 => data <= "10010101";
        when 681 => data <= "10000100";
        when 682 => data <= "00000001";
        when 683 => data <= "00101101";
        when 684 => data <= "01011001";
        when 685 => data <= "00010010";
        when 686 => data <= "10100100";
        when 687 => data <= "10010101";
        when 688 => data <= "01010101";
        when 689 => data <= "01001110";
        when 690 => data <= "01010010";
        when 691 => data <= "00100101";
        when 692 => data <= "01000101";
        when 693 => data <= "00011001";
        when 694 => data <= "01010010";
        when 695 => data <= "01010001";
        when 696 => data <= "01010101";
        when 697 => data <= "01000101";
        when 698 => data <= "00010011";
        when 699 => data <= "01010000";
        when 700 => data <= "11010001";
        when 701 => data <= "01110101";
        when 702 => data <= "00001101";
        when 703 => data <= "00100010";
        when 704 => data <= "01010110";
        when 705 => data <= "00010111";
        when 706 => data <= "11111100";
        when 707 => data <= "00001001";
        when 708 => data <= "01111011";
        when 709 => data <= "01001110";
        when 710 => data <= "11010000";
        when 711 => data <= "00100100";
        when 712 => data <= "01101101";
        when 713 => data <= "01001011";
        when 714 => data <= "01001110";
        when 715 => data <= "11010101";
        when 716 => data <= "00110100";
        when 717 => data <= "00001001";
        when 718 => data <= "00100010";
        when 719 => data <= "01001111";
        when 720 => data <= "00110010";
        when 721 => data <= "11100100";
        when 722 => data <= "00001111";
        when 723 => data <= "01011000";
        when 724 => data <= "01011111";
        when 725 => data <= "11110011";
        when 726 => data <= "01000100";
        when 727 => data <= "11001011";
        when 728 => data <= "00100011";
        when 729 => data <= "11000110";
        when 730 => data <= "10010100";
        when 731 => data <= "00001100";
        when 732 => data <= "11101011";
        when 733 => data <= "00110010";
        when 734 => data <= "01000010";
        when 735 => data <= "10010001";
        when 736 => data <= "00001100";
        when 737 => data <= "10100001";
        when 738 => data <= "01100111";
        when 739 => data <= "11010000";
        when 740 => data <= "01010010";
        when 741 => data <= "11101100";
        when 742 => data <= "11010001";
        when 743 => data <= "00001110";
        when 744 => data <= "01000111";
        when 745 => data <= "11010011";
        when 746 => data <= "11001101";
        when 747 => data <= "11000001";
        when 748 => data <= "00101110";
        when 749 => data <= "11011111";
        when 750 => data <= "01010011";
        when 751 => data <= "01100100";
        when 752 => data <= "11110001";
        when 753 => data <= "00111111";
        when 754 => data <= "11010110";
        when 755 => data <= "01010000";
        when 756 => data <= "11101101";
        when 757 => data <= "00111101";
        when 758 => data <= "00011001";
        when 759 => data <= "01010001";
        when 760 => data <= "00010000";
        when 761 => data <= "00011101";
        when 762 => data <= "01001001";
        when 763 => data <= "00001001";
        when 764 => data <= "01000000";
        when 765 => data <= "11010010";
        when 766 => data <= "10001100";
        when 767 => data <= "10101111";
        when 768 => data <= "01101111";
        when 769 => data <= "11001010";
        when 770 => data <= "01110010";
        when 771 => data <= "11100100";
        when 772 => data <= "11000111";
        when 773 => data <= "00011011";
        when 774 => data <= "11011110";
        when 775 => data <= "01110111";
        when 776 => data <= "01111100";
        when 777 => data <= "11001101";
        when 778 => data <= "00001111";
        when 779 => data <= "11010001";
        when 780 => data <= "11110110";
        when 781 => data <= "01010101";
        when 782 => data <= "00010011";
        when 783 => data <= "01011111";
        when 784 => data <= "01010101";
        when 785 => data <= "01110110";
        when 786 => data <= "11010101";
        when 787 => data <= "11010111";
        when 788 => data <= "00010101";
        when 789 => data <= "11000111";
        when 790 => data <= "11010000";
        when 791 => data <= "10001101";
        when 792 => data <= "10100111";
        when 793 => data <= "01011001";
        when 794 => data <= "11000011";
        when 795 => data <= "11010101";
        when 796 => data <= "01001101";
        when 797 => data <= "11101001";
        when 798 => data <= "01111101";
        when 799 => data <= "11000101";
        when 800 => data <= "10011111";
        when 801 => data <= "11111111";
        when 802 => data <= "11111111";
        when 803 => data <= "11111111";
        when 804 => data <= "11111111";
        when 805 => data <= "11111111";
        when 806 => data <= "11111111";
        when 807 => data <= "11111111";
        when 808 => data <= "11111111";
        when 809 => data <= "11111111";
        when 810 => data <= "11111111";
        when 811 => data <= "11111111";
        when 812 => data <= "11111111";
        when 813 => data <= "11111111";
        when 814 => data <= "11111111";
        when 815 => data <= "11111111";
        when 816 => data <= "11111111";
        when 817 => data <= "11111111";
        when 818 => data <= "11111111";
        when 819 => data <= "11111111";
        when 820 => data <= "11111111";
        when 821 => data <= "11111111";
        when 822 => data <= "11111111";
        when 823 => data <= "11111111";
        when 824 => data <= "11111111";
        when 825 => data <= "11111111";
        when 826 => data <= "11111111";
        when 827 => data <= "11111111";
        when 828 => data <= "11111111";
        when 829 => data <= "11111111";
        when 830 => data <= "11111111";
        when 831 => data <= "11111111";
        when 832 => data <= "11111111";
        when 833 => data <= "11111111";
        when 834 => data <= "11111111";
        when 835 => data <= "11111111";
        when 836 => data <= "11111111";
        when 837 => data <= "11111111";
        when 838 => data <= "11111111";
        when 839 => data <= "11111111";
        when 840 => data <= "11111111";
        when 841 => data <= "11111111";
        when 842 => data <= "11111111";
        when 843 => data <= "11111111";
        when 844 => data <= "11111111";
        when 845 => data <= "11111111";
        when 846 => data <= "11111111";
        when 847 => data <= "11111111";
        when 848 => data <= "11111111";
        when 849 => data <= "11111111";
        when 850 => data <= "11111111";
        when 851 => data <= "11111111";
        when 852 => data <= "11111111";
        when 853 => data <= "11111111";
        when 854 => data <= "11111111";
        when 855 => data <= "11111111";
        when 856 => data <= "11111111";
        when 857 => data <= "11111111";
        when 858 => data <= "11111111";
        when 859 => data <= "11111111";
        when 860 => data <= "11111111";
        when 861 => data <= "11111111";
        when 862 => data <= "11111111";
        when 863 => data <= "11111111";
        when 864 => data <= "11111111";
        when 865 => data <= "11111111";
        when 866 => data <= "11111111";
        when 867 => data <= "11111111";
        when 868 => data <= "11111111";
        when 869 => data <= "11111111";
        when 870 => data <= "11111111";
        when 871 => data <= "11111111";
        when 872 => data <= "11111111";
        when 873 => data <= "11111111";
        when 874 => data <= "11111111";
        when 875 => data <= "11111111";
        when 876 => data <= "11111111";
        when 877 => data <= "11111111";
        when 878 => data <= "11111111";
        when 879 => data <= "11111111";
        when 880 => data <= "11111111";
        when 881 => data <= "11111111";
        when 882 => data <= "11111111";
        when 883 => data <= "11111111";
        when 884 => data <= "11111111";
        when 885 => data <= "11111111";
        when 886 => data <= "11111111";
        when 887 => data <= "11111111";
        when 888 => data <= "11111111";
        when 889 => data <= "11111111";
        when 890 => data <= "11111111";
        when 891 => data <= "11111111";
        when 892 => data <= "11111111";
        when 893 => data <= "11111111";
        when 894 => data <= "11111111";
        when 895 => data <= "11111111";
        when 896 => data <= "11111111";
        when 897 => data <= "11111111";
        when 898 => data <= "11111111";
        when 899 => data <= "11111111";
        when 900 => data <= "11111111";
        when 901 => data <= "11111111";
        when 902 => data <= "11111111";
        when 903 => data <= "11111111";
        when 904 => data <= "11111111";
        when 905 => data <= "11111111";
        when 906 => data <= "11111111";
        when 907 => data <= "11111111";
        when 908 => data <= "11111111";
        when 909 => data <= "11111111";
        when 910 => data <= "11111111";
        when 911 => data <= "11111111";
        when 912 => data <= "11111111";
        when 913 => data <= "11111111";
        when 914 => data <= "11111111";
        when 915 => data <= "11111111";
        when 916 => data <= "11111111";
        when 917 => data <= "11111111";
        when 918 => data <= "11111111";
        when 919 => data <= "11111111";
        when 920 => data <= "11111111";
        when 921 => data <= "11111111";
        when 922 => data <= "11111111";
        when 923 => data <= "11111111";
        when 924 => data <= "11111111";
        when 925 => data <= "11111111";
        when 926 => data <= "11111111";
        when 927 => data <= "11111111";
        when 928 => data <= "11111111";
        when 929 => data <= "11111111";
        when 930 => data <= "11111111";
        when 931 => data <= "11111111";
        when 932 => data <= "11111111";
        when 933 => data <= "11111111";
        when 934 => data <= "11111111";
        when 935 => data <= "11111111";
        when 936 => data <= "11111111";
        when 937 => data <= "11111111";
        when 938 => data <= "11111111";
        when 939 => data <= "11111111";
        when 940 => data <= "11111111";
        when 941 => data <= "11111111";
        when 942 => data <= "11111111";
        when 943 => data <= "11111111";
        when 944 => data <= "11111111";
        when 945 => data <= "11111111";
        when 946 => data <= "11111111";
        when 947 => data <= "11111111";
        when 948 => data <= "11111111";
        when 949 => data <= "11111111";
        when 950 => data <= "11111111";
        when 951 => data <= "11111111";
        when 952 => data <= "11111111";
        when 953 => data <= "11111111";
        when 954 => data <= "11111111";
        when 955 => data <= "11111111";
        when 956 => data <= "11111111";
        when 957 => data <= "11111111";
        when 958 => data <= "11111111";
        when 959 => data <= "11111111";
        when 960 => data <= "11111111";
        when 961 => data <= "11111111";
        when 962 => data <= "11111111";
        when 963 => data <= "11111111";
        when 964 => data <= "11111111";
        when 965 => data <= "11111111";
        when 966 => data <= "11111111";
        when 967 => data <= "11111111";
        when 968 => data <= "11111111";
        when 969 => data <= "11111111";
        when 970 => data <= "11111111";
        when 971 => data <= "11111111";
        when 972 => data <= "11111111";
        when 973 => data <= "11111111";
        when 974 => data <= "11111111";
        when 975 => data <= "11111111";
        when 976 => data <= "11111111";
        when 977 => data <= "11111111";
        when 978 => data <= "11111111";
        when 979 => data <= "11111111";
        when 980 => data <= "11111111";
        when 981 => data <= "11111111";
        when 982 => data <= "11111111";
        when 983 => data <= "11111111";
        when 984 => data <= "11111111";
        when 985 => data <= "11111111";
        when 986 => data <= "11111111";
        when 987 => data <= "11111111";
        when 988 => data <= "11111111";
        when 989 => data <= "11111111";
        when 990 => data <= "11111111";
        when 991 => data <= "11111111";
        when 992 => data <= "11111111";
        when 993 => data <= "11111111";
        when 994 => data <= "11111111";
        when 995 => data <= "11111111";
        when 996 => data <= "11111111";
        when 997 => data <= "11111111";
        when 998 => data <= "11111111";
        when 999 => data <= "11111111";
        when 1000 => data <= "11111111";
        when 1001 => data <= "11111111";
        when 1002 => data <= "11111111";
        when 1003 => data <= "11111111";
        when 1004 => data <= "11111111";
        when 1005 => data <= "11111111";
        when 1006 => data <= "11111111";
        when 1007 => data <= "11111111";
        when 1008 => data <= "11111111";
        when 1009 => data <= "11111111";
        when 1010 => data <= "11111111";
        when 1011 => data <= "11111111";
        when 1012 => data <= "11111111";
        when 1013 => data <= "11111111";
        when 1014 => data <= "11111111";
        when 1015 => data <= "11111111";
        when 1016 => data <= "11111111";
        when 1017 => data <= "11111111";
        when 1018 => data <= "11111111";
        when 1019 => data <= "11111111";
        when 1020 => data <= "11111111";
        when 1021 => data <= "11111111";
        when 1022 => data <= "11111111";
        when 1023 => data <= "11111111";
        when 1024 => data <= "11111111";
        when 1025 => data <= "11111111";
        when 1026 => data <= "11111111";
        when 1027 => data <= "11111111";
        when 1028 => data <= "11111111";
        when 1029 => data <= "11111111";
        when 1030 => data <= "11111111";
        when 1031 => data <= "11111111";
        when 1032 => data <= "11111111";
        when 1033 => data <= "11111111";
        when 1034 => data <= "11111111";
        when 1035 => data <= "11111111";
        when 1036 => data <= "11111111";
        when 1037 => data <= "11111111";
        when 1038 => data <= "11111111";
        when 1039 => data <= "11111111";
        when 1040 => data <= "11111111";
        when 1041 => data <= "11111111";
        when 1042 => data <= "11111111";
        when 1043 => data <= "11111111";
        when 1044 => data <= "11111111";
        when 1045 => data <= "11111111";
        when 1046 => data <= "11111111";
        when 1047 => data <= "11111111";
        when 1048 => data <= "11111111";
        when 1049 => data <= "11111111";
        when 1050 => data <= "11111111";
        when 1051 => data <= "11111111";
        when 1052 => data <= "11111111";
        when 1053 => data <= "11111111";
        when 1054 => data <= "11111111";
        when 1055 => data <= "11111111";
        when 1056 => data <= "11111111";
        when 1057 => data <= "11111111";
        when 1058 => data <= "11111111";
        when 1059 => data <= "11111111";
        when 1060 => data <= "11111111";
        when 1061 => data <= "11111111";
        when 1062 => data <= "11111111";
        when 1063 => data <= "11111111";
        when 1064 => data <= "11111111";
        when 1065 => data <= "11111111";
        when 1066 => data <= "11111111";
        when 1067 => data <= "11111111";
        when 1068 => data <= "11111111";
        when 1069 => data <= "11111111";
        when 1070 => data <= "11111111";
        when 1071 => data <= "11111111";
        when 1072 => data <= "11111111";
        when 1073 => data <= "11111111";
        when 1074 => data <= "11111111";
        when 1075 => data <= "11111111";
        when 1076 => data <= "11111111";
        when 1077 => data <= "11111111";
        when 1078 => data <= "11111111";
        when 1079 => data <= "11111111";
        when 1080 => data <= "11111111";
        when 1081 => data <= "11111111";
        when 1082 => data <= "11111111";
        when 1083 => data <= "11111111";
        when 1084 => data <= "11111111";
        when 1085 => data <= "11111111";
        when 1086 => data <= "11111111";
        when 1087 => data <= "11111111";
        when 1088 => data <= "11111111";
        when 1089 => data <= "11111111";
        when 1090 => data <= "11111111";
        when 1091 => data <= "11111111";
        when 1092 => data <= "11111111";
        when 1093 => data <= "11111111";
        when 1094 => data <= "11111111";
        when 1095 => data <= "11111111";
        when 1096 => data <= "11111111";
        when 1097 => data <= "11111111";
        when 1098 => data <= "11111111";
        when 1099 => data <= "11111111";
        when 1100 => data <= "11111110";
        when 1101 => data <= "00000000";
        when 1102 => data <= "00000000";
        when 1103 => data <= "00000000";
        when 1104 => data <= "00000000";
        when 1105 => data <= "00000000";
        when 1106 => data <= "00000000";
        when 1107 => data <= "00000000";
        when 1108 => data <= "00000000";
        when 1109 => data <= "00000000";
        when 1110 => data <= "00000000";
        when 1111 => data <= "00000000";
        when 1112 => data <= "00000000";
        when 1113 => data <= "00000000";
        when 1114 => data <= "00000000";
        when 1115 => data <= "00000000";
        when 1116 => data <= "00000000";
        when 1117 => data <= "00000000";
        when 1118 => data <= "00000000";
        when 1119 => data <= "00000000";
        when 1120 => data <= "00000000";
        when 1121 => data <= "00000000";
        when 1122 => data <= "00000000";
        when 1123 => data <= "00000000";
        when 1124 => data <= "00000000";
        when 1125 => data <= "00000000";
        when 1126 => data <= "00000000";
        when 1127 => data <= "00000000";
        when 1128 => data <= "00000000";
        when 1129 => data <= "00000000";
        when 1130 => data <= "00000000";
        when 1131 => data <= "00000000";
        when 1132 => data <= "00000000";
        when 1133 => data <= "00000000";
        when 1134 => data <= "00000000";
        when 1135 => data <= "00000000";
        when 1136 => data <= "00000000";
        when 1137 => data <= "00000000";
        when 1138 => data <= "00000000";
        when 1139 => data <= "00000000";
        when 1140 => data <= "00000000";
        when 1141 => data <= "00000000";
        when 1142 => data <= "00000000";
        when 1143 => data <= "00000000";
        when 1144 => data <= "00000000";
        when 1145 => data <= "00000000";
        when 1146 => data <= "00000000";
        when 1147 => data <= "00000000";
        when 1148 => data <= "00000000";
        when 1149 => data <= "00000000";
        when 1150 => data <= "00000000";
        when 1151 => data <= "00000000";
        when 1152 => data <= "00000000";
        when 1153 => data <= "00000000";
        when 1154 => data <= "00000000";
        when 1155 => data <= "00000000";
        when 1156 => data <= "00000000";
        when 1157 => data <= "00000000";
        when 1158 => data <= "00000000";
        when 1159 => data <= "00000000";
        when 1160 => data <= "00000000";
        when 1161 => data <= "00000000";
        when 1162 => data <= "00000000";
        when 1163 => data <= "00000000";
        when 1164 => data <= "00000000";
        when 1165 => data <= "00000000";
        when 1166 => data <= "00000000";
        when 1167 => data <= "00000000";
        when 1168 => data <= "00000000";
        when 1169 => data <= "00000000";
        when 1170 => data <= "00000000";
        when 1171 => data <= "00000000";
        when 1172 => data <= "00000000";
        when 1173 => data <= "00000000";
        when 1174 => data <= "00000000";
        when 1175 => data <= "00000000";
        when 1176 => data <= "00000000";
        when 1177 => data <= "00000000";
        when 1178 => data <= "00000000";
        when 1179 => data <= "00000000";
        when 1180 => data <= "00000000";
        when 1181 => data <= "00000000";
        when 1182 => data <= "00000000";
        when 1183 => data <= "00000000";
        when 1184 => data <= "00000000";
        when 1185 => data <= "00000000";
        when 1186 => data <= "00000000";
        when 1187 => data <= "00000000";
        when 1188 => data <= "00000000";
        when 1189 => data <= "00000000";
        when 1190 => data <= "00000000";
        when 1191 => data <= "00000000";
        when 1192 => data <= "00000000";
        when 1193 => data <= "00000000";
        when 1194 => data <= "00000000";
        when 1195 => data <= "00000000";
        when 1196 => data <= "00000000";
        when 1197 => data <= "00000000";
        when 1198 => data <= "00000000";
        when 1199 => data <= "00000000";
        when 1200 => data <= "00000000";
        when 1201 => data <= "00000000";
        when 1202 => data <= "00000000";
        when 1203 => data <= "00000000";
        when 1204 => data <= "00000000";
        when 1205 => data <= "00000000";
        when 1206 => data <= "00000000";
        when 1207 => data <= "00000000";
        when 1208 => data <= "00000000";
        when 1209 => data <= "00000000";
        when 1210 => data <= "00000000";
        when 1211 => data <= "00000000";
        when 1212 => data <= "00000000";
        when 1213 => data <= "00000000";
        when 1214 => data <= "00000000";
        when 1215 => data <= "00000000";
        when 1216 => data <= "00000000";
        when 1217 => data <= "00000000";
        when 1218 => data <= "00000000";
        when 1219 => data <= "00000000";
        when 1220 => data <= "00000000";
        when 1221 => data <= "00000000";
        when 1222 => data <= "00000000";
        when 1223 => data <= "00000000";
        when 1224 => data <= "00000000";
        when 1225 => data <= "00000000";
        when 1226 => data <= "00000000";
        when 1227 => data <= "00000000";
        when 1228 => data <= "00000000";
        when 1229 => data <= "00000000";
        when 1230 => data <= "00000000";
        when 1231 => data <= "00000000";
        when 1232 => data <= "00000000";
        when 1233 => data <= "00000000";
        when 1234 => data <= "00000000";
        when 1235 => data <= "00000000";
        when 1236 => data <= "00000000";
        when 1237 => data <= "00000000";
        when 1238 => data <= "00000000";
        when 1239 => data <= "00000000";
        when 1240 => data <= "00000000";
        when 1241 => data <= "00000000";
        when 1242 => data <= "00000000";
        when 1243 => data <= "00000000";
        when 1244 => data <= "00000000";
        when 1245 => data <= "00000000";
        when 1246 => data <= "00000000";
        when 1247 => data <= "00000000";
        when 1248 => data <= "00000000";
        when 1249 => data <= "00000000";
        when 1250 => data <= "00000000";
        when 1251 => data <= "00000000";
        when 1252 => data <= "00000000";
        when 1253 => data <= "00000000";
        when 1254 => data <= "00000000";
        when 1255 => data <= "00000000";
        when 1256 => data <= "00000000";
        when 1257 => data <= "00000000";
        when 1258 => data <= "00000000";
        when 1259 => data <= "00000000";
        when 1260 => data <= "00000000";
        when 1261 => data <= "00000000";
        when 1262 => data <= "00000000";
        when 1263 => data <= "00000000";
        when 1264 => data <= "00000000";
        when 1265 => data <= "00000000";
        when 1266 => data <= "00000000";
        when 1267 => data <= "00000000";
        when 1268 => data <= "00000000";
        when 1269 => data <= "00000000";
        when 1270 => data <= "00000000";
        when 1271 => data <= "00000000";
        when 1272 => data <= "00000000";
        when 1273 => data <= "00000000";
        when 1274 => data <= "00000000";
        when 1275 => data <= "00000000";
        when 1276 => data <= "00000000";
        when 1277 => data <= "00000000";
        when 1278 => data <= "00000000";
        when 1279 => data <= "00000000";
        when 1280 => data <= "00000000";
        when 1281 => data <= "00000000";
        when 1282 => data <= "00000000";
        when 1283 => data <= "00000000";
        when 1284 => data <= "00000000";
        when 1285 => data <= "00000000";
        when 1286 => data <= "00000000";
        when 1287 => data <= "00000000";
        when 1288 => data <= "00000000";
        when 1289 => data <= "00000000";
        when 1290 => data <= "00000000";
        when 1291 => data <= "00000000";
        when 1292 => data <= "00000000";
        when 1293 => data <= "00000000";
        when 1294 => data <= "00000000";
        when 1295 => data <= "00000000";
        when 1296 => data <= "00000000";
        when 1297 => data <= "00000000";
        when 1298 => data <= "00000000";
        when 1299 => data <= "00000000";
        when 1300 => data <= "00000000";
        when 1301 => data <= "00000000";
        when 1302 => data <= "00000000";
        when 1303 => data <= "00000000";
        when 1304 => data <= "00000000";
        when 1305 => data <= "00000000";
        when 1306 => data <= "00000000";
        when 1307 => data <= "00000000";
        when 1308 => data <= "00000000";
        when 1309 => data <= "00000000";
        when 1310 => data <= "00000000";
        when 1311 => data <= "00000000";
        when 1312 => data <= "00000000";
        when 1313 => data <= "00000000";
        when 1314 => data <= "00000000";
        when 1315 => data <= "00000000";
        when 1316 => data <= "00000000";
        when 1317 => data <= "00000000";
        when 1318 => data <= "00000000";
        when 1319 => data <= "00000000";
        when 1320 => data <= "00000000";
        when 1321 => data <= "00000000";
        when 1322 => data <= "00000000";
        when 1323 => data <= "00000000";
        when 1324 => data <= "00000000";
        when 1325 => data <= "00000000";
        when 1326 => data <= "00000000";
        when 1327 => data <= "00000000";
        when 1328 => data <= "00000000";
        when 1329 => data <= "00000000";
        when 1330 => data <= "00000000";
        when 1331 => data <= "00000000";
        when 1332 => data <= "00000000";
        when 1333 => data <= "00000000";
        when 1334 => data <= "00000000";
        when 1335 => data <= "00000000";
        when 1336 => data <= "00000000";
        when 1337 => data <= "00000000";
        when 1338 => data <= "00000000";
        when 1339 => data <= "00000000";
        when 1340 => data <= "00000000";
        when 1341 => data <= "00000000";
        when 1342 => data <= "00000000";
        when 1343 => data <= "00000000";
        when 1344 => data <= "00000000";
        when 1345 => data <= "00000000";
        when 1346 => data <= "00000000";
        when 1347 => data <= "00000000";
        when 1348 => data <= "00000000";
        when 1349 => data <= "00000000";
        when 1350 => data <= "00000000";
        when 1351 => data <= "00000000";
        when 1352 => data <= "00000000";
        when 1353 => data <= "00000000";
        when 1354 => data <= "00000000";
        when 1355 => data <= "00000000";
        when 1356 => data <= "00000000";
        when 1357 => data <= "00000000";
        when 1358 => data <= "00000000";
        when 1359 => data <= "00000000";
        when 1360 => data <= "00000000";
        when 1361 => data <= "00000000";
        when 1362 => data <= "00000000";
        when 1363 => data <= "00000000";
        when 1364 => data <= "00000000";
        when 1365 => data <= "00000000";
        when 1366 => data <= "00000000";
        when 1367 => data <= "00000000";
        when 1368 => data <= "00000000";
        when 1369 => data <= "00000000";
        when 1370 => data <= "00000000";
        when 1371 => data <= "00000000";
        when 1372 => data <= "00000000";
        when 1373 => data <= "00000000";
        when 1374 => data <= "00000000";
        when 1375 => data <= "00000000";
        when 1376 => data <= "00000000";
        when 1377 => data <= "00000000";
        when 1378 => data <= "00000000";
        when 1379 => data <= "00000000";
        when 1380 => data <= "00000000";
        when 1381 => data <= "00000000";
        when 1382 => data <= "00000000";
        when 1383 => data <= "00000000";
        when 1384 => data <= "00000000";
        when 1385 => data <= "00000000";
        when 1386 => data <= "00000000";
        when 1387 => data <= "00000000";
        when 1388 => data <= "00000000";
        when 1389 => data <= "00000000";
        when 1390 => data <= "00000000";
        when 1391 => data <= "00000000";
        when 1392 => data <= "00000000";
        when 1393 => data <= "00000000";
        when 1394 => data <= "00000000";
        when 1395 => data <= "00000000";
        when 1396 => data <= "00000000";
        when 1397 => data <= "00000000";
        when 1398 => data <= "00000000";
        when 1399 => data <= "00000000";
        when 1400 => data <= "00000000";
        when 1401 => data <= "00111111";
        when 1402 => data <= "11111111";
        when 1403 => data <= "11111111";
        when 1404 => data <= "11111111";
        when 1405 => data <= "11111111";
        when 1406 => data <= "11111111";
        when 1407 => data <= "11111111";
        when 1408 => data <= "11111111";
        when 1409 => data <= "11111111";
        when 1410 => data <= "11111111";
        when 1411 => data <= "11111111";
        when 1412 => data <= "11111111";
        when 1413 => data <= "11111111";
        when 1414 => data <= "11111111";
        when 1415 => data <= "11111111";
        when 1416 => data <= "11111111";
        when 1417 => data <= "11111111";
        when 1418 => data <= "11111111";
        when 1419 => data <= "11111111";
        when 1420 => data <= "11111111";
        when 1421 => data <= "11111111";
        when 1422 => data <= "11111111";
        when 1423 => data <= "11111111";
        when 1424 => data <= "11111111";
        when 1425 => data <= "11111111";
        when 1426 => data <= "11111111";
        when 1427 => data <= "11111111";
        when 1428 => data <= "11111111";
        when 1429 => data <= "11111111";
        when 1430 => data <= "11111111";
        when 1431 => data <= "11111111";
        when 1432 => data <= "11111111";
        when 1433 => data <= "11111111";
        when 1434 => data <= "11111111";
        when 1435 => data <= "11111111";
        when 1436 => data <= "11111111";
        when 1437 => data <= "11111111";
        when 1438 => data <= "11111111";
        when 1439 => data <= "11111111";
        when 1440 => data <= "11111111";
        when 1441 => data <= "11111111";
        when 1442 => data <= "11111111";
        when 1443 => data <= "11111111";
        when 1444 => data <= "11111111";
        when 1445 => data <= "11111111";
        when 1446 => data <= "11111111";
        when 1447 => data <= "11111111";
        when 1448 => data <= "11111111";
        when 1449 => data <= "11111111";
        when 1450 => data <= "11111111";
        when 1451 => data <= "11111111";
        when 1452 => data <= "11111111";
        when 1453 => data <= "11111111";
        when 1454 => data <= "11111111";
        when 1455 => data <= "11111111";
        when 1456 => data <= "11111111";
        when 1457 => data <= "11111111";
        when 1458 => data <= "11111111";
        when 1459 => data <= "11111111";
        when 1460 => data <= "11111111";
        when 1461 => data <= "11111111";
        when 1462 => data <= "11111111";
        when 1463 => data <= "11111111";
        when 1464 => data <= "11111111";
        when 1465 => data <= "11111111";
        when 1466 => data <= "11111111";
        when 1467 => data <= "11111111";
        when 1468 => data <= "11111111";
        when 1469 => data <= "11111111";
        when 1470 => data <= "11111111";
        when 1471 => data <= "11111111";
        when 1472 => data <= "11111111";
        when 1473 => data <= "11111111";
        when 1474 => data <= "11111111";
        when 1475 => data <= "11111111";
        when 1476 => data <= "11111111";
        when 1477 => data <= "11111111";
        when 1478 => data <= "11111111";
        when 1479 => data <= "11111111";
        when 1480 => data <= "11111111";
        when 1481 => data <= "11111111";
        when 1482 => data <= "11111111";
        when 1483 => data <= "11111111";
        when 1484 => data <= "11111111";
        when 1485 => data <= "11111111";
        when 1486 => data <= "11111111";
        when 1487 => data <= "11111111";
        when 1488 => data <= "11111111";
        when 1489 => data <= "11111111";
        when 1490 => data <= "11111111";
        when 1491 => data <= "11111111";
        when 1492 => data <= "11111111";
        when 1493 => data <= "11111111";
        when 1494 => data <= "11111111";
        when 1495 => data <= "11111111";
        when 1496 => data <= "11111111";
        when 1497 => data <= "11111111";
        when 1498 => data <= "11111111";
        when 1499 => data <= "11111111";
        when 1500 => data <= "11111111";
        when 1501 => data <= "11111111";
        when 1502 => data <= "11111111";
        when 1503 => data <= "11111111";
        when 1504 => data <= "11111111";
        when 1505 => data <= "11111111";
        when 1506 => data <= "11111111";
        when 1507 => data <= "11111111";
        when 1508 => data <= "11111111";
        when 1509 => data <= "11111111";
        when 1510 => data <= "11111111";
        when 1511 => data <= "11111111";
        when 1512 => data <= "11111111";
        when 1513 => data <= "11111111";
        when 1514 => data <= "11111111";
        when 1515 => data <= "11111111";
        when 1516 => data <= "11111111";
        when 1517 => data <= "11111111";
        when 1518 => data <= "11111111";
        when 1519 => data <= "11111111";
        when 1520 => data <= "11111111";
        when 1521 => data <= "11111111";
        when 1522 => data <= "11111111";
        when 1523 => data <= "11111111";
        when 1524 => data <= "11111111";
        when 1525 => data <= "11111111";
        when 1526 => data <= "11111111";
        when 1527 => data <= "11111111";
        when 1528 => data <= "11111111";
        when 1529 => data <= "11111111";
        when 1530 => data <= "11111111";
        when 1531 => data <= "11111111";
        when 1532 => data <= "11111111";
        when 1533 => data <= "11111111";
        when 1534 => data <= "11111111";
        when 1535 => data <= "11111111";
        when 1536 => data <= "11111111";
        when 1537 => data <= "11111111";
        when 1538 => data <= "11111111";
        when 1539 => data <= "11111111";
        when 1540 => data <= "11111111";
        when 1541 => data <= "11111111";
        when 1542 => data <= "11111111";
        when 1543 => data <= "11111111";
        when 1544 => data <= "11111111";
        when 1545 => data <= "11111111";
        when 1546 => data <= "11111111";
        when 1547 => data <= "11111111";
        when 1548 => data <= "11111111";
        when 1549 => data <= "11111111";
        when 1550 => data <= "11111111";
        when 1551 => data <= "11111111";
        when 1552 => data <= "11111111";
        when 1553 => data <= "11111111";
        when 1554 => data <= "11111111";
        when 1555 => data <= "11111111";
        when 1556 => data <= "11111111";
        when 1557 => data <= "11111111";
        when 1558 => data <= "11111111";
        when 1559 => data <= "11111111";
        when 1560 => data <= "11111111";
        when 1561 => data <= "11111111";
        when 1562 => data <= "11111111";
        when 1563 => data <= "11111111";
        when 1564 => data <= "11111111";
        when 1565 => data <= "11111111";
        when 1566 => data <= "11111111";
        when 1567 => data <= "11111111";
        when 1568 => data <= "11111111";
        when 1569 => data <= "11111111";
        when 1570 => data <= "11111111";
        when 1571 => data <= "11111111";
        when 1572 => data <= "11111111";
        when 1573 => data <= "11111111";
        when 1574 => data <= "11111111";
        when 1575 => data <= "11111111";
        when 1576 => data <= "11111111";
        when 1577 => data <= "11111111";
        when 1578 => data <= "11111111";
        when 1579 => data <= "11111111";
        when 1580 => data <= "11111111";
        when 1581 => data <= "11111111";
        when 1582 => data <= "11111111";
        when 1583 => data <= "11111111";
        when 1584 => data <= "11111111";
        when 1585 => data <= "11111111";
        when 1586 => data <= "11111111";
        when 1587 => data <= "11111111";
        when 1588 => data <= "11111111";
        when 1589 => data <= "11111111";
        when 1590 => data <= "11111111";
        when 1591 => data <= "11111111";
        when 1592 => data <= "11111111";
        when 1593 => data <= "11111111";
        when 1594 => data <= "11111111";
        when 1595 => data <= "11111111";
        when 1596 => data <= "11111111";
        when 1597 => data <= "11111111";
        when 1598 => data <= "11111111";
        when 1599 => data <= "11111111";
        when 1600 => data <= "11111111";
        when 1601 => data <= "11111111";
        when 1602 => data <= "11111111";
        when 1603 => data <= "11111111";
        when 1604 => data <= "11111111";
        when 1605 => data <= "11111111";
        when 1606 => data <= "11111111";
        when 1607 => data <= "11111111";
        when 1608 => data <= "11111111";
        when 1609 => data <= "11111111";
        when 1610 => data <= "11111111";
        when 1611 => data <= "11111111";
        when 1612 => data <= "11111111";
        when 1613 => data <= "11111111";
        when 1614 => data <= "11111111";
        when 1615 => data <= "11111111";
        when 1616 => data <= "11111111";
        when 1617 => data <= "11111111";
        when 1618 => data <= "11111111";
        when 1619 => data <= "11111111";
        when 1620 => data <= "11111111";
        when 1621 => data <= "11111111";
        when 1622 => data <= "11111111";
        when 1623 => data <= "11111111";
        when 1624 => data <= "11111111";
        when 1625 => data <= "11111111";
        when 1626 => data <= "11110001";
        when 1627 => data <= "11011111";
        when 1628 => data <= "11111111";
        when 1629 => data <= "11111111";
        when 1630 => data <= "11111111";
        when 1631 => data <= "11111111";
        when 1632 => data <= "11111111";
        when 1633 => data <= "11111111";
        when 1634 => data <= "11111111";
        when 1635 => data <= "11111111";
        when 1636 => data <= "11111111";
        when 1637 => data <= "11111111";
        when 1638 => data <= "11111111";
        when 1639 => data <= "11111111";
        when 1640 => data <= "11111111";
        when 1641 => data <= "11111111";
        when 1642 => data <= "11111111";
        when 1643 => data <= "11111111";
        when 1644 => data <= "11111111";
        when 1645 => data <= "11111111";
        when 1646 => data <= "11111111";
        when 1647 => data <= "11111111";
        when 1648 => data <= "11111111";
        when 1649 => data <= "11111111";
        when 1650 => data <= "11111111";
        when 1651 => data <= "11111111";
        when 1652 => data <= "11111111";
        when 1653 => data <= "11111111";
        when 1654 => data <= "11111111";
        when 1655 => data <= "11111111";
        when 1656 => data <= "11111111";
        when 1657 => data <= "11111111";
        when 1658 => data <= "11111111";
        when 1659 => data <= "11111111";
        when 1660 => data <= "11111111";
        when 1661 => data <= "11111111";
        when 1662 => data <= "11111111";
        when 1663 => data <= "11111111";
        when 1664 => data <= "11111111";
        when 1665 => data <= "11111111";
        when 1666 => data <= "11111111";
        when 1667 => data <= "11111111";
        when 1668 => data <= "11111111";
        when 1669 => data <= "11111111";
        when 1670 => data <= "11111111";
        when 1671 => data <= "11111111";
        when 1672 => data <= "11111111";
        when 1673 => data <= "11111111";
        when 1674 => data <= "11111111";
        when 1675 => data <= "11111111";
        when 1676 => data <= "11111111";
        when 1677 => data <= "11111111";
        when 1678 => data <= "11111111";
        when 1679 => data <= "11111111";
        when 1680 => data <= "11111111";
        when 1681 => data <= "11111111";
        when 1682 => data <= "11111111";
        when 1683 => data <= "11111111";
        when 1684 => data <= "11111111";
        when 1685 => data <= "11111111";
        when 1686 => data <= "11111111";
        when 1687 => data <= "11111111";
        when 1688 => data <= "11111111";
        when 1689 => data <= "11111111";
        when 1690 => data <= "11111111";
        when 1691 => data <= "11111111";
        when 1692 => data <= "11111111";
        when 1693 => data <= "11111111";
        when 1694 => data <= "11111111";
        when 1695 => data <= "11111111";
        when 1696 => data <= "11111111";
        when 1697 => data <= "11111111";
        when 1698 => data <= "11111111";
        when 1699 => data <= "11111111";
        when 1700 => data <= "11111111";
        when 1701 => data <= "11111111";
        when 1702 => data <= "11111111";
        when 1703 => data <= "11111111";
        when 1704 => data <= "11111111";
        when 1705 => data <= "11111111";
        when 1706 => data <= "11111111";
        when 1707 => data <= "11111111";
        when 1708 => data <= "11111111";
        when 1709 => data <= "11111111";
        when 1710 => data <= "11111111";
        when 1711 => data <= "11111111";
        when 1712 => data <= "11111111";
        when 1713 => data <= "11111111";
        when 1714 => data <= "11111111";
        when 1715 => data <= "11111111";
        when 1716 => data <= "11111111";
        when 1717 => data <= "11111111";
        when 1718 => data <= "11111111";
        when 1719 => data <= "11111111";
        when 1720 => data <= "11111111";
        when 1721 => data <= "11111111";
        when 1722 => data <= "11111111";
        when 1723 => data <= "11111111";
        when 1724 => data <= "11111111";
        when 1725 => data <= "11111111";
        when 1726 => data <= "11111111";
        when 1727 => data <= "11111111";
        when 1728 => data <= "11111111";
        when 1729 => data <= "11111111";
        when 1730 => data <= "11111111";
        when 1731 => data <= "11111111";
        when 1732 => data <= "11111111";
        when 1733 => data <= "11111111";
        when 1734 => data <= "11111111";
        when 1735 => data <= "11111111";
        when 1736 => data <= "11111111";
        when 1737 => data <= "11111111";
        when 1738 => data <= "11111111";
        when 1739 => data <= "11111111";
        when 1740 => data <= "11111111";
        when 1741 => data <= "11111111";
        when 1742 => data <= "11111111";
        when 1743 => data <= "11111111";
        when 1744 => data <= "11111111";
        when 1745 => data <= "11111111";
        when 1746 => data <= "11111111";
        when 1747 => data <= "11111111";
        when 1748 => data <= "11111111";
        when 1749 => data <= "11111111";
        when 1750 => data <= "11111111";
        when 1751 => data <= "11111111";
        when 1752 => data <= "11111111";
        when 1753 => data <= "11111111";
        when 1754 => data <= "11111111";
        when 1755 => data <= "11111111";
        when 1756 => data <= "11111111";
        when 1757 => data <= "11111111";
        when 1758 => data <= "11111111";
        when 1759 => data <= "11111111";
        when 1760 => data <= "11111111";
        when 1761 => data <= "11111111";
        when 1762 => data <= "11111111";
        when 1763 => data <= "11111111";
        when 1764 => data <= "11111111";
        when 1765 => data <= "11111111";
        when 1766 => data <= "11111111";
        when 1767 => data <= "11111111";
        when 1768 => data <= "11111111";
        when 1769 => data <= "11111111";
        when 1770 => data <= "11111111";
        when 1771 => data <= "11111111";
        when 1772 => data <= "11111111";
        when 1773 => data <= "11111111";
        when 1774 => data <= "11111111";
        when 1775 => data <= "11111111";
        when 1776 => data <= "11111111";
        when 1777 => data <= "11111111";
        when 1778 => data <= "11111111";
        when 1779 => data <= "11111111";
        when 1780 => data <= "11111111";
        when 1781 => data <= "11111111";
        when 1782 => data <= "11111111";
        when 1783 => data <= "11111111";
        when 1784 => data <= "11111111";
        when 1785 => data <= "11111111";
        when 1786 => data <= "11111111";
        when 1787 => data <= "11111111";
        when 1788 => data <= "11111111";
        when 1789 => data <= "11111111";
        when 1790 => data <= "11111111";
        when 1791 => data <= "11111111";
        when 1792 => data <= "11111111";
        when 1793 => data <= "11111111";
        when 1794 => data <= "11111111";
        when 1795 => data <= "11111111";
        when 1796 => data <= "11111111";
        when 1797 => data <= "11111111";
        when 1798 => data <= "11111111";
        when 1799 => data <= "11111111";
        when 1800 => data <= "11111111";
        when 1801 => data <= "11111111";
        when 1802 => data <= "11111111";
        when 1803 => data <= "11111111";
        when 1804 => data <= "11111111";
        when 1805 => data <= "11111111";
        when 1806 => data <= "11111111";
        when 1807 => data <= "11111111";
        when 1808 => data <= "11111111";
        when 1809 => data <= "11111111";
        when 1810 => data <= "11111111";
        when 1811 => data <= "11111111";
        when 1812 => data <= "11111111";
        when 1813 => data <= "11111111";
        when 1814 => data <= "11111111";
        when 1815 => data <= "11111111";
        when 1816 => data <= "11111111";
        when 1817 => data <= "11111111";
        when 1818 => data <= "11111111";
        when 1819 => data <= "11111111";
        when 1820 => data <= "11111111";
        when 1821 => data <= "11111111";
        when 1822 => data <= "11111111";
        when 1823 => data <= "11111111";
        when 1824 => data <= "11111111";
        when 1825 => data <= "11111111";
        when 1826 => data <= "11111111";
        when 1827 => data <= "11111111";
        when 1828 => data <= "11111111";
        when 1829 => data <= "11111111";
        when 1830 => data <= "11111111";
        when 1831 => data <= "11111111";
        when 1832 => data <= "11111111";
        when 1833 => data <= "11111111";
        when 1834 => data <= "11111111";
        when 1835 => data <= "11111111";
        when 1836 => data <= "11111111";
        when 1837 => data <= "11111111";
        when 1838 => data <= "11111111";
        when 1839 => data <= "11111111";
        when 1840 => data <= "11111111";
        when 1841 => data <= "11111111";
        when 1842 => data <= "11111111";
        when 1843 => data <= "11111111";
        when 1844 => data <= "11111111";
        when 1845 => data <= "11111111";
        when 1846 => data <= "11111111";
        when 1847 => data <= "11111111";
        when 1848 => data <= "11111111";
        when 1849 => data <= "11111111";
        when 1850 => data <= "11111111";
        when 1851 => data <= "11111111";
        when 1852 => data <= "11111111";
        when 1853 => data <= "00101010";
        when 1854 => data <= "01010100";
        when 1855 => data <= "01010001";
        when 1856 => data <= "10010101";
        when 1857 => data <= "00100101";
        when 1858 => data <= "00010101";
        when 1859 => data <= "01010100";
        when 1860 => data <= "01010001";
        when 1861 => data <= "00110101";
        when 1862 => data <= "00001101";
        when 1863 => data <= "00010111";
        when 1864 => data <= "01010000";
        when 1865 => data <= "11010000";
        when 1866 => data <= "00000100";
        when 1867 => data <= "00000001";
        when 1868 => data <= "00111000";
        when 1869 => data <= "01011111";
        when 1870 => data <= "11110111";
        when 1871 => data <= "11111100";
        when 1872 => data <= "00000001";
        when 1873 => data <= "00011100";
        when 1874 => data <= "01011111";
        when 1875 => data <= "11110111";
        when 1876 => data <= "11111100";
        when 1877 => data <= "00000001";
        when 1878 => data <= "00000000";
        when 1879 => data <= "01000000";
        when 1880 => data <= "00010100";
        when 1881 => data <= "00000101";
        when 1882 => data <= "00000001";
        when 1883 => data <= "00000000";
        when 1884 => data <= "01000000";
        when 1885 => data <= "00010000";
        when 1886 => data <= "00000100";
        when 1887 => data <= "00000001";
        when 1888 => data <= "01101100";
        when 1889 => data <= "01000101";
        when 1890 => data <= "11010001";
        when 1891 => data <= "11110100";
        when 1892 => data <= "00000001";
        when 1893 => data <= "01111001";
        when 1894 => data <= "01000101";
        when 1895 => data <= "00110001";
        when 1896 => data <= "01001101";
        when 1897 => data <= "10111111";
        when 1898 => data <= "00100010";
        when 1899 => data <= "01001110";
        when 1900 => data <= "01010001";
        when 1901 => data <= "00010101";
        when 1902 => data <= "00101001";
        when 1903 => data <= "01001111";
        when 1904 => data <= "11000011";
        when 1905 => data <= "10010100";
        when 1906 => data <= "11100101";
        when 1907 => data <= "10101001";
        when 1908 => data <= "00100101";
        when 1909 => data <= "11000011";
        when 1910 => data <= "00010001";
        when 1911 => data <= "00110100";
        when 1912 => data <= "10000001";
        when 1913 => data <= "01111110";
        when 1914 => data <= "11000000";
        when 1915 => data <= "10010110";
        when 1916 => data <= "10010100";
        when 1917 => data <= "00000001";
        when 1918 => data <= "00010001";
        when 1919 => data <= "01010000";
        when 1920 => data <= "00110111";
        when 1921 => data <= "01111101";
        when 1922 => data <= "11110001";
        when 1923 => data <= "00110100";
        when 1924 => data <= "01000011";
        when 1925 => data <= "01110111";
        when 1926 => data <= "11000100";
        when 1927 => data <= "00000101";
        when 1928 => data <= "01111010";
        when 1929 => data <= "01010011";
        when 1930 => data <= "10010001";
        when 1931 => data <= "01010100";
        when 1932 => data <= "10011001";
        when 1933 => data <= "00101101";
        when 1934 => data <= "11001000";
        when 1935 => data <= "00010001";
        when 1936 => data <= "10110100";
        when 1937 => data <= "11111101";
        when 1938 => data <= "01011000";
        when 1939 => data <= "01010001";
        when 1940 => data <= "01010111";
        when 1941 => data <= "11111101";
        when 1942 => data <= "11011101";
        when 1943 => data <= "01011100";
        when 1944 => data <= "01000001";
        when 1945 => data <= "11010111";
        when 1946 => data <= "01110100";
        when 1947 => data <= "00101101";
        when 1948 => data <= "00110001";
        when 1949 => data <= "11000110";
        when 1950 => data <= "10110111";
        when 1951 => data <= "00001101";
        when 1952 => data <= "00000011";
        when 1953 => data <= "00000101";
        when 1954 => data <= "11011110";
        when 1955 => data <= "11110110";
        when 1956 => data <= "10100100";
        when 1957 => data <= "10001101";
        when 1958 => data <= "01101000";
        when 1959 => data <= "01010101";
        when 1960 => data <= "11010100";
        when 1961 => data <= "11100100";
        when 1962 => data <= "00110111";
        when 1963 => data <= "01011100";
        when 1964 => data <= "11010100";
        when 1965 => data <= "10010000";
        when 1966 => data <= "11110101";
        when 1967 => data <= "01110001";
        when 1968 => data <= "00001111";
        when 1969 => data <= "01001000";
        when 1970 => data <= "11110001";
        when 1971 => data <= "01000101";
        when 1972 => data <= "11010001";
        when 1973 => data <= "00011110";
        when 1974 => data <= "11011100";
        when 1975 => data <= "10010111";
        when 1976 => data <= "00100100";
        when 1977 => data <= "00111101";
        when 1978 => data <= "01010011";
        when 1979 => data <= "01000110";
        when 1980 => data <= "01110101";
        when 1981 => data <= "11011100";
        when 1982 => data <= "01111111";
        when 1983 => data <= "01011010";
        when 1984 => data <= "11010101";
        when 1985 => data <= "01110010";
        when 1986 => data <= "10010100";
        when 1987 => data <= "10011001";
        when 1988 => data <= "00000101";
        when 1989 => data <= "11001110";
        when 1990 => data <= "10110000";
        when 1991 => data <= "11101100";
        when 1992 => data <= "01100011";
        when 1993 => data <= "01001011";
        when 1994 => data <= "11011010";
        when 1995 => data <= "01110110";
        when 1996 => data <= "10001101";
        when 1997 => data <= "00011011";
        when 1998 => data <= "00001101";
        when 1999 => data <= "11001101";
        when 2000 => data <= "10010111";
        when 2001 => data <= "10110100";
        when 2002 => data <= "00111101";
        when 2003 => data <= "01101000";
        when 2004 => data <= "11000001";
        when 2005 => data <= "00010011";
        when 2006 => data <= "10001100";
        when 2007 => data <= "00000111";
        when 2008 => data <= "00110100";
        when 2009 => data <= "11000010";
        when 2010 => data <= "00110101";
        when 2011 => data <= "10001101";
        when 2012 => data <= "01011101";
        when 2013 => data <= "00001011";
        when 2014 => data <= "01011010";
        when 2015 => data <= "11110011";
        when 2016 => data <= "01110101";
        when 2017 => data <= "00000001";
        when 2018 => data <= "01011000";
        when 2019 => data <= "11011111";
        when 2020 => data <= "10110010";
        when 2021 => data <= "11101101";
        when 2022 => data <= "00110001";
        when 2023 => data <= "00101000";
        when 2024 => data <= "11010100";
        when 2025 => data <= "00110101";
        when 2026 => data <= "10001101";
        when 2027 => data <= "00111011";
        when 2028 => data <= "01101010";
        when 2029 => data <= "11010110";
        when 2030 => data <= "11110000";
        when 2031 => data <= "10110100";
        when 2032 => data <= "00111101";
        when 2033 => data <= "01011000";
        when 2034 => data <= "11001000";
        when 2035 => data <= "11010001";
        when 2036 => data <= "00110101";
        when 2037 => data <= "11110111";
        when 2038 => data <= "01110000";
        when 2039 => data <= "01001100";
        when 2040 => data <= "10010000";
        when 2041 => data <= "10001101";
        when 2042 => data <= "11000111";
        when 2043 => data <= "00110111";
        when 2044 => data <= "01001000";
        when 2045 => data <= "11110100";
        when 2046 => data <= "01001100";
        when 2047 => data <= "01100001";
        when 2048 => data <= "00011000";
        when 2049 => data <= "01010010";
        when 2050 => data <= "10010001";
        when 2051 => data <= "10101101";
        when 2052 => data <= "00100111";
        when 2053 => data <= "01111111";
        when 2054 => data <= "11011111";
        when 2055 => data <= "10010011";
        when 2056 => data <= "11001100";
        when 2057 => data <= "00110011";
        when 2058 => data <= "01011000";
        when 2059 => data <= "11000001";
        when 2060 => data <= "11110001";
        when 2061 => data <= "10110100";
        when 2062 => data <= "11101001";
        when 2063 => data <= "00010001";
        when 2064 => data <= "11001111";
        when 2065 => data <= "00110110";
        when 2066 => data <= "11010100";
        when 2067 => data <= "00010111";
        when 2068 => data <= "01010000";
        when 2069 => data <= "01010001";
        when 2070 => data <= "10010001";
        when 2071 => data <= "11010101";
        when 2072 => data <= "01001011";
        when 2073 => data <= "01001111";
        when 2074 => data <= "11000000";
        when 2075 => data <= "01110110";
        when 2076 => data <= "00110100";
        when 2077 => data <= "01111111";
        when 2078 => data <= "01001111";
        when 2079 => data <= "01010000";
        when 2080 => data <= "11110010";
        when 2081 => data <= "00111100";
        when 2082 => data <= "00101111";
        when 2083 => data <= "00101011";
        when 2084 => data <= "11001000";
        when 2085 => data <= "01110111";
        when 2086 => data <= "01101100";
        when 2087 => data <= "00000111";
        when 2088 => data <= "00101111";
        when 2089 => data <= "01000000";
        when 2090 => data <= "10010001";
        when 2091 => data <= "01001101";
        when 2092 => data <= "01000101";
        when 2093 => data <= "01000101";
        when 2094 => data <= "11010100";
        when 2095 => data <= "01010110";
        when 2096 => data <= "11000101";
        when 2097 => data <= "10011111";
        when 2098 => data <= "01100010";
        when 2099 => data <= "01010101";
        when 2100 => data <= "00110011";
        when 2101 => data <= "10101101";
        when 2102 => data <= "11100111";
        when 2103 => data <= "00000100";
        when 2104 => data <= "11000001";
        when 2105 => data <= "01010001";
        when 2106 => data <= "00100100";
        when 2107 => data <= "11011101";
        when 2108 => data <= "01111101";
        when 2109 => data <= "01000001";
        when 2110 => data <= "01110100";
        when 2111 => data <= "00111100";
        when 2112 => data <= "00110111";
        when 2113 => data <= "01101100";
        when 2114 => data <= "11010100";
        when 2115 => data <= "01110011";
        when 2116 => data <= "01110100";
        when 2117 => data <= "00000101";
        when 2118 => data <= "00001110";
        when 2119 => data <= "01000111";
        when 2120 => data <= "00010010";
        when 2121 => data <= "10101101";
        when 2122 => data <= "00111001";
        when 2123 => data <= "00100101";
        when 2124 => data <= "11011111";
        when 2125 => data <= "10110000";
        when 2126 => data <= "00101100";
        when 2127 => data <= "01010011";
        when 2128 => data <= "00110101";
        when 2129 => data <= "01001011";
        when 2130 => data <= "00110111";
        when 2131 => data <= "00010100";
        when 2132 => data <= "10101011";
        when 2133 => data <= "01011011";
        when 2134 => data <= "01001110";
        when 2135 => data <= "01110111";
        when 2136 => data <= "10110100";
        when 2137 => data <= "01110011";
        when 2138 => data <= "01010010";
        when 2139 => data <= "01011111";
        when 2140 => data <= "10110100";
        when 2141 => data <= "10101100";
        when 2142 => data <= "10100011";
        when 2143 => data <= "00001101";
        when 2144 => data <= "11011001";
        when 2145 => data <= "11110110";
        when 2146 => data <= "01001101";
        when 2147 => data <= "11111001";
        when 2148 => data <= "01111011";
        when 2149 => data <= "01011010";
        when 2150 => data <= "01110010";
        when 2151 => data <= "10000101";
        when 2152 => data <= "00001011";
        when 2153 => data <= "00000000";
        when 2154 => data <= "01000001";
        when 2155 => data <= "01110001";
        when 2156 => data <= "01001100";
        when 2157 => data <= "10110011";
        when 2158 => data <= "01100000";
        when 2159 => data <= "11000111";
        when 2160 => data <= "11110111";
        when 2161 => data <= "10110100";
        when 2162 => data <= "11000011";
        when 2163 => data <= "00010000";
        when 2164 => data <= "11011010";
        when 2165 => data <= "10110100";
        when 2166 => data <= "00010100";
        when 2167 => data <= "00011101";
        when 2168 => data <= "00010000";
        when 2169 => data <= "01011000";
        when 2170 => data <= "00010110";
        when 2171 => data <= "01010101";
        when 2172 => data <= "10001001";
        when 2173 => data <= "01111011";
        when 2174 => data <= "01001101";
        when 2175 => data <= "00110001";
        when 2176 => data <= "10110100";
        when 2177 => data <= "10001101";
        when 2178 => data <= "01110110";
        when 2179 => data <= "11010101";
        when 2180 => data <= "00010101";
        when 2181 => data <= "10000100";
        when 2182 => data <= "11000111";
        when 2183 => data <= "01100111";
        when 2184 => data <= "01000110";
        when 2185 => data <= "01010111";
        when 2186 => data <= "11100100";
        when 2187 => data <= "01101101";
        when 2188 => data <= "01000010";
        when 2189 => data <= "11001100";
        when 2190 => data <= "11010000";
        when 2191 => data <= "01111101";
        when 2192 => data <= "01110011";
        when 2193 => data <= "00101001";
        when 2194 => data <= "11011101";
        when 2195 => data <= "11010110";
        when 2196 => data <= "00011100";
        when 2197 => data <= "01011111";
        when 2198 => data <= "01001111";
        when 2199 => data <= "01010101";
        when 2200 => data <= "10010010";
        when 2201 => data <= "11001100";
        when 2202 => data <= "11001011";
        when 2203 => data <= "00110010";
        when 2204 => data <= "11001011";
        when 2205 => data <= "10110100";
        when 2206 => data <= "00100101";
        when 2207 => data <= "10010111";
        when 2208 => data <= "01111101";
        when 2209 => data <= "11011000";
        when 2210 => data <= "01110001";
        when 2211 => data <= "11101100";
        when 2212 => data <= "00000111";
        when 2213 => data <= "11111111";
        when 2214 => data <= "11111111";
        when 2215 => data <= "11111111";
        when 2216 => data <= "11111111";
        when 2217 => data <= "11111111";
        when 2218 => data <= "11111111";
        when 2219 => data <= "11111111";
        when 2220 => data <= "11111111";
        when 2221 => data <= "11111111";
        when 2222 => data <= "11111111";
        when 2223 => data <= "11111111";
        when 2224 => data <= "11111111";
        when 2225 => data <= "11111111";
        when 2226 => data <= "11111111";
        when 2227 => data <= "11111111";
        when 2228 => data <= "11111111";
        when 2229 => data <= "11111111";
        when 2230 => data <= "11111111";
        when 2231 => data <= "11111111";
        when 2232 => data <= "11111111";
        when 2233 => data <= "11111111";
        when 2234 => data <= "11111111";
        when 2235 => data <= "11111111";
        when 2236 => data <= "11111111";
        when 2237 => data <= "11111111";
        when 2238 => data <= "11111111";
        when 2239 => data <= "11111111";
        when 2240 => data <= "11111111";
        when 2241 => data <= "11111111";
        when 2242 => data <= "11111111";
        when 2243 => data <= "11111111";
        when 2244 => data <= "11111111";
        when 2245 => data <= "11111111";
        when 2246 => data <= "11111111";
        when 2247 => data <= "11111111";
        when 2248 => data <= "11111111";
        when 2249 => data <= "11111111";
        when 2250 => data <= "11111111";
        when 2251 => data <= "11111111";
        when 2252 => data <= "11111111";
        when 2253 => data <= "11111111";
        when 2254 => data <= "11111111";
        when 2255 => data <= "11111111";
        when 2256 => data <= "11111111";
        when 2257 => data <= "11111111";
        when 2258 => data <= "11111111";
        when others => data <= "00000000";
      end case;
    
    end if; -- rising_edge

  end process;


  --
  -- FILEIO
  --
  -- u_FileIO_FCh : entity work.Replay_FileIO_FCh_Generic
  -- port map (
  --   -- clocks
  --   i_clk                 => i_clk_sys,
  --   i_ena                 => i_ena_sys,
  --   i_rst                 => i_rst_sys,

  --   -- FileIO / Syscon interface
  --   i_fch_to_core         => i_fch_to_core,
  --   o_fch_fm_core         => o_fch_fm_core,

  --   -- to user space
  --   i_req                 => fileio_req,
  --   o_ack_req             => fileio_ack_req,
  --   o_ack_trans           => fileio_ack_trans, -- transfer done
  --   o_trans_err           => fileio_trans_err, -- aborted, truncated, seek error

  --   -- below latched on ack
  --   i_dir                 => '0', -- read only
  --   i_chan                => "00",
  --   i_addr                => fileio_addr,
  --   i_size                => fileio_size,
  --   o_size0               => fileio_src_size,

  --   -- Reading
  --   i_fifo_to_core_flush  => '0',
  --   o_fifo_to_core_data   => fileio_data,
  --   i_fifo_to_core_taken  => fileio_taken,
  --   o_fifo_to_core_valid  => fileio_valid,
  --   o_fifo_to_core_level  => fileio_rx_level,
  --   o_fifo_to_core_overfl => fileio_rx_overfl,

  --   -- Writing
  --   i_fifo_fm_core_flush  => '0',
  --   i_fifo_fm_core_data   => (others => '0'),
  --   i_fifo_fm_core_we     => '0',
  --   o_fifo_fm_core_level  => open
  --   );
  
  -- -- request size is 512 16 bits words
  -- fileio_size <= x"0400";

  -- -- Enable/pause data request via the Generic FileIO entity
  -- p_fileio_req : process(i_clk_sys, i_rst_sys)
  -- begin   
  --   if (i_rst_sys = '1') then
  --     fileio_addr <= (others => '0');
  --     fileio_req  <= '0';
  --     fileio_req_state <= S_IDLE;
  --   elsif rising_edge(i_clk_sys) then
  --     if (i_ena_sys = '1') then
  --       fileio_req  <= '0';

  --       if (i_fcha_cfg.inserted(0) = '0') then
  --         fileio_addr <= (others => '0');
  --         fileio_req_state <= S_IDLE;
  --       else
  --         case fileio_req_state is
  --           when S_IDLE =>
  --             if (fileio_rx_level(9) = '0') then -- <hf
  --               fileio_req  <= '1'; -- note, request only sent when ack received
  --             end if;
  --             if (fileio_ack_req = '1') then
  --               fileio_req_state <= S_WAIT;
  --             end if;

  --           when S_WAIT =>
  --             if (fileio_ack_trans = '1') then
  --               if (red_or(fileio_trans_err) = '1') then
  --                 fileio_addr <= (others => '0');
  --               else
  --                 fileio_addr <= fileio_addr + fileio_size;
  --               end if;
  --               fileio_req_state <= S_IDLE;
  --             end if;

  --           when others => null;
  --         end case;
  --       end if;
  --     end if;
  --   end if;
  -- end process;

  -- -- Transfer available sample data from FIFO out to audio subsystem  
  -- p_fileio_reader : process(i_clk_sys, i_rst_sys)
  -- begin
  --   if (i_rst_sys = '1') then
  --           fileio_sample_cnt <= "00";
  --           fileio_taken      <= '0';
  --           sample_audio_l   <= (others => '0');
  --           sample_audio_r   <= (others => '0');
  --   elsif rising_edge(i_clk_sys) then


  --     if (i_ena_sys = '1') then
        
  --       sys_audio_taken_sync_old <= sys_audio_taken_sync;
  --       sys_audio_taken_sync <= audio_taken_sync;
        
  --       fileio_taken <= '0';
  --       case fileio_sample_cnt is
  --         when "00" =>
  --           if (fileio_valid = '1') then
  --             fileio_taken <= '1';
  --             sample_audio_l   <= fileio_data( 7 downto 0) & fileio_data(15 downto 8) & x"00";
  --             --o_audio_l  <= fileio_data(15 downto 0)  & x"00";
  --             fileio_sample_cnt <= "01";
  --           end if;
  --         when "01" => -- wait for taken to update valid
  --             fileio_sample_cnt <= "10";

  --         when "10" =>
  --           if (fileio_valid = '1') then
  --             fileio_taken <= '1';
  --             sample_audio_r   <= fileio_data( 7 downto 0) & fileio_data(15 downto 8) & x"00";
  --             --o_audio_r   <= fileio_data(15 downto 0) & x"00";
  --             fileio_sample_cnt <= "11";
  --           end if;
  --         when "11" => -- ready
  --           if (sys_audio_taken_sync /= sys_audio_taken_sync_old) then              
              
  --             fileio_sample_cnt <= "00";
  --           end if;
  --         when others => null;
  --       end case;
  --     end if;
  --   end if;

  -- end process;
    
  -- p_audio_out : process
  -- begin    
  --   wait until rising_edge(i_clk_aud);

  --   if (i_ena_aud = '1') then
  --     o_audio_l <= sample_audio_l;
  --     o_audio_r <= sample_audio_r;

  --     -- Stretch taken pulse to sync with reader process
  --     if (i_audio_taken = '1') then
  --       audio_taken_sync <= not audio_taken_sync;
  --     end if;
  --   end if;

  -- end process;

end RTL;