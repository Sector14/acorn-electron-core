-- Acorn Electron ULA
-- Ferranti 12C021 Custom

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

  use work.Replay_Pack.all;
  use work.Replay_VideoTiming_Pack.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ULA_12C021 is
  port (
    foo : out bit1
  );
end;

architecture RTL of ULA_12C021 is
begin


-- RAM

-- 
end;
